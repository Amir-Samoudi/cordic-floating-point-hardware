library verilog;
use verilog.vl_types.all;
entity TB_reciprocal is
end TB_reciprocal;
