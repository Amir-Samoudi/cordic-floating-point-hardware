library verilog;
use verilog.vl_types.all;
entity TB_square_root_float is
end TB_square_root_float;
