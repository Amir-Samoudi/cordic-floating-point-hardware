library verilog;
use verilog.vl_types.all;
entity TB_reciprocal_float is
end TB_reciprocal_float;
