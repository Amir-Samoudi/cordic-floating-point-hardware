library verilog;
use verilog.vl_types.all;
entity TB_cordic_linear is
end TB_cordic_linear;
